--nao faz nada